----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 2019/11/11 15:31:13
-- Design Name: 
-- Module Name: Imem - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Imem is
 Port (
        PCin: in std_logic_vector(31 downto 0);
        rst: in std_logic;
        clk: in std_logic;
        addressout: out std_logic_vector(31 downto 0);
        ishalt: out std_logic
  );
end Imem;

architecture Behavioral of Imem is

TYPE rom IS ARRAY (0 TO 895) OF STD_LOGIC_VECTOR(7 DOWNTO 0); 
--CONSTANT irom: rom:=rom'( "00010000","00000001","00000000","01111011","00010000","00000010","00000001","11001000");
CONSTANT irom: rom:=rom'("11111100","00000000","00000000","00000000","00011100","00000001","00000000","00110100","00011100","00000010","00000000","00110101","00000000","00100000","00001001","11010101","00000000","00100000","00001001","11010101","00000000","00100010","00001000","10010101","00011100","00000010","00000000","00110110","00011100","00000011","00000000","00110111","00000000","01000000","00010001","11010101","00000000","01000000","00010001","11010101","00000000","01000011","00010000","10010101","00011100","00011101","00000000","00000000","00011100","00011110","00000000","00011010","00000011","10100000","11101001","11010101","00000011","10100000","11101001","11010101","00000011","10111110","11101000","10010101","00011100","00011110","00000000","00000001","00011100","00011111","00000000","00011011","00000011","11000000","11110001","11010101","00000011","11000000","11110001","11010101","00000011","11011111","11110000","10010101","00000000","00111101","00001000","00010101","00000000","01011110","00010000","00010101","00010000","00000011","00000000","00000001","00010000","00011111","00000000","00000001","00010000","00000100","00000000","00011001","00000000","01111111","00011000","00010101","00011100","01100101","00000000","00000000","00011100","01100110","00000000","00011010","00000000","10100000","00101001","11010101","00000000","10100000","00101001","11010101","00000000","10100110","00101000","10010101","00001100","01000111","00000000","00011111","00000000","00000000","01000000","00010101","00101000","11101000","00000000","00111110","00000001","00011111","01000000","00010101","00101000","11101000","00000000","00111110","00000001","00011111","01000000","00010101","00101000","11101000","00000000","00111110","00000001","00011111","01000000","00010101","00101000","11101000","00000000","00111110","00000001","00011111","01000000","00010101","00101000","11101000","00000000","00111110","00000001","00011111","01000000","00010101","00101000","11101000","00000000","00111110","00000001","00011111","01000000","00010101","00101000","11101000","00000000","00111110","00000001","00011111","01000000","00010101","00101000","11101000","00000000","00111110","00000001","00011111","01000000","00010101","00101000","11101000","00000000","00111110","00000001","00011111","01000000","00010101","00101000","11101000","00000000","00111111","00000001","00011111","01000000","00010101","00101000","11101000","00000000","01000000","00000001","00011111","01000000","00010101","00101000","11101000","00000000","01000001","00000001","00011111","01000000","00010101","00101000","11101000","00000000","01000010","00000001","00011111","01000000","00010101","00101000","11101000","00000000","01000011","00000001","00011111","01000000","00010101","00101000","11101000","00000000","01000100","00000001","00011111","01000000","00010101","00101000","11101000","00000000","01000101","00000001","00011111","01000000","00010101","00101000","11101000","00000000","01000111","00000001","00011111","01000000","00010101","00101000","11101000","00000000","01001001","00000001","00011111","01000000","00010101","00101000","11101000","00000000","01001011","00000001","00011111","01000000","00010101","00101000","11101000","00000000","01001101","00000001","00011111","01000000","00010101","00101000","11101000","00000000","01001111","00000001","00011111","01000000","00010101","00101000","11101000","00000000","01010001","00000001","00011111","01000000","00010101","00101000","11101000","00000000","01010011","00000001","00011111","01000000","00010101","00101000","11101000","00000000","01010110","00000001","00011111","01000000","00010101","00101000","11101000","00000000","01011001","00000001","00011111","01000000","00010101","00101000","11101000","00000000","01011100","00000001","00011111","01000000","00010101","00101000","11101000","00000000","01011111","00000001","00011111","01000000","00010101","00101000","11101000","00000000","01100010","00000001","00011111","01000000","00010101","00101000","11101000","00000000","01100101","00000001","00011111","01000000","00010101","00101000","11101000","00000000","01101000","00000001","00011111","01000000","00010101","00101000","11101000","00000000","01101100","00000001","00011111","01000000","00010101","00101000","11101000","00000000","01110000","00000000","00100010","00001000","00010000","00110000","00000000","00000000","01110100","00000000","00100010","00001000","01010000","00110000","00000000","00000000","01110010","00000000","00100010","00001000","10010000","00110000","00000000","00000000","01110000","00000000","00100010","00001000","11010000","00110000","00000000","00000000","01101110","00000000","00100010","00001001","00010000","00110000","00000000","00000000","01101100","00000000","00100010","00001001","01010000","00110000","00000000","00000000","01101010","00000000","00100010","00001001","10010000","00110000","00000000","00000000","01101000","00000000","00100010","00001001","11010000","00110000","00000000","00000000","01100110","00000000","00100010","00001001","11010000","00000000","00100000","00001000","01010101","00110000","00000000","00000000","01100011","00000000","00100010","00001001","11010000","00000000","00100000","00001000","10010101","00110000","00000000","00000000","01100000","00000000","00100010","00001001","11010000","00000000","00100000","00001000","11010101","00110000","00000000","00000000","01011101","00000000","00100010","00001001","11010000","00000000","00100000","00001001","00010101","00110000","00000000","00000000","01011010","00000000","00100010","00001001","11010000","00000000","00100000","00001001","01010101","00110000","00000000","00000000","01010111","00000000","00100010","00001001","11010000","00000000","00100000","00001001","10010101","00110000","00000000","00000000","01010100","00000000","00100010","00001001","11010000","00000000","00100000","00001001","11010101","00110000","00000000","00000000","01010001","00000000","00100010","00001001","11010000","00000000","00100000","00001001","11010101","00000000","00100000","00001000","01010101","00110000","00000000","00000000","01001101","00000000","00100010","00001001","11010000","00000000","00100000","00001001","11010101","00000000","00100000","00001000","10010101","00110000","00000000","00000000","01001001","00000000","00100010","00001001","11010000","00000000","00100000","00001001","11010101","00000000","00100000","00001000","11010101","00110000","00000000","00000000","01000101","00000000","00100010","00001001","11010000","00000000","00100000","00001001","11010101","00000000","00100000","00001001","00010101","00110000","00000000","00000000","01000001","00000000","00100010","00001001","11010000","00000000","00100000","00001001","11010101","00000000","00100000","00001001","01010101","00110000","00000000","00000000","00111101","00000000","00100010","00001001","11010000","00000000","00100000","00001001","11010101","00000000","00100000","00001001","10010101","00110000","00000000","00000000","00111001","00000000","00100010","00001001","11010000","00000000","00100000","00001001","11010101","00000000","00100000","00001001","11010101","00110000","00000000","00000000","00110101","00000000","00100010","00001001","11010000","00000000","00100000","00001001","11010101","00000000","00100000","00001001","11010101","00000000","00100000","00001000","01010101","00110000","00000000","00000000","00110000","00000000","00100010","00001001","11010000","00000000","00100000","00001001","11010101","00000000","00100000","00001001","11010101","00000000","00100000","00001000","10010101","00110000","00000000","00000000","00101011","00000000","00100010","00001001","11010000","00000000","00100000","00001001","11010101","00000000","00100000","00001001","11010101","00000000","00100000","00001000","11010101","00110000","00000000","00000000","00100110","00000000","00100010","00001001","11010000","00000000","00100000","00001001","11010101","00000000","00100000","00001001","11010101","00000000","00100000","00001001","00010101","00110000","00000000","00000000","00100001","00000000","00100010","00001001","11010000","00000000","00100000","00001001","11010101","00000000","00100000","00001001","11010101","00000000","00100000","00001001","01010101","00110000","00000000","00000000","00011100","00000000","00100010","00001001","11010000","00000000","00100000","00001001","11010101","00000000","00100000","00001001","11010101","00000000","00100000","00001001","10010101","00110000","00000000","00000000","00010111","00000000","00100010","00001001","11010000","00000000","00100000","00001001","11010101","00000000","00100000","00001001","11010101","00000000","00100000","00001001","11010101","00110000","00000000","00000000","00010010","00000000","00100010","00001001","11010000","00000000","00100000","00001001","11010101","00000000","00100000","00001001","11010101","00000000","00100000","00001001","11010101","00000000","00100000","00001000","01010101","00110000","00000000","00000000","00001100","00000000","00100010","00001001","11010000","00000000","00100000","00001001","11010101","00000000","00100000","00001001","11010101","00000000","00100000","00001001","11010101","00000000","00100000","00001000","10010101","00110000","00000000","00000000","00000110","00000000","00100010","00001001","11010000","00000000","00100000","00001001","11010101","00000000","00100000","00001001","11010101","00000000","00100000","00001001","11010101","00000000","00100000","00001000","11010101","00110000","00000000","00000000","00000000","00000000","00100101","00001000","00010101","00000000","00100000","01001000","00010101","00000000","01000000","00001000","00010101","00000001","00100000","00010000","00010101","00101100","01100100","11111111","00111110","00000000","00100000","01011001","11010101","00000001","01100000","01011001","11010101","00000001","01100010","01011000","10010101","11111100","00000000","00000000","00000000"
);
--signal count:std_logic_vector(2 downto 0);
signal count:std_logic_vector(31 downto 0):=x"00000000";
signal address_judge:std_logic_vector(31 downto 0);

begin
count<=PCin;
--address_judge<=irom(CONV_INTEGER(count))& irom(CONV_INTEGER(count+'1'))& irom(CONV_INTEGER(count+"10")) & irom(CONV_INTEGER(count+"11"));
ishalt<='1' when address_judge="11111100000000000000000000000000"            else '0';
address_judge<=irom(CONV_INTEGER(count))& irom(CONV_INTEGER(count+'1'))& irom(CONV_INTEGER(count+"10")) & irom(CONV_INTEGER(count+"11"));
addressout<=address_judge;
--process(clk,rst)
--begin
--    if(clk' event and clk='1')then
    --address_judge<=irom(CONV_INTEGER(count)/4);
       
--    end if;
--end process;
    --addressout<=address_judge;
--    if (rst = '1') then
--        addressout <="00000000000000000000000000000000";
--        ishalt<='0';
--        --count<=0;
--    --elsif(clk 'event and clk='1') then
--        --if(count="11111100000000000000000000000000");
--    elsif (address_judge="11111100000000000000000000000000")then 
--        ishalt<='1';
--    else
--        address_judge<=irom(CONV_INTEGER(count))& irom(CONV_INTEGER(count+'1'))& irom(CONV_INTEGER(count+"10")) & irom(CONV_INTEGER(count+"11"));
--        addressout<=address_judge;
--    end if;
--end process;



end Behavioral;